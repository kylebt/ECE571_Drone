module rpmctrl(clk, resetn, angle, alt_rpm, rpm_set);
input clk, resetn;
input [15:0] angle, alt_rpm;
output [15:0] rpm_set;

// multiply alt_rpm by angle
endmodule