module dirctrl(clk, resetn, cmds, angle);
input clk, resetn;
input [2:0] cmds;
output [15:0];

// based on cmds output angle value
endmodule

