module altctrl(clk, resetn, altcmd, alt_rpm);
input clk, resetn;
input [2:0] altcmd;
output [15:0] alt_rpm;

// see notes on DroneController module drawing
endmodule